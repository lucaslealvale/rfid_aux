
module RFID_NIOS (
	clk_clk,
	reset_reset_n,
	rfid_tx_rfid);	

	input		clk_clk;
	input		reset_reset_n;
	output		rfid_tx_rfid;
endmodule
